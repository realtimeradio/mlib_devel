`timescale 1ns/100ps

module htg_ad9213_quad_top #(
  parameter USE_FMC_A=1'b1,
  parameter USE_FMC_B=1'b1,
  parameter USE_FMC_C=1'b1,
  parameter USE_FMC_D=1'b0
  ) (
  // 200MHz external clock
  input         clk_200_p,
  input         clk_200_n,
  // Software reset, driven from Simulink
  input         reset,
  // External UART pins -- always on FMC C
  input         uart_txd,
  output        uart_rxd,
  //// FMC A
  // HMC
  output        hmc_a_sync,
  output        hmc_a_reset,
  inout         hmc_a_gpio1,
  inout         hmc_a_gpio2,
  inout         hmc_a_gpio3,
  inout         hmc_a_gpio4,
  // SPI
  output        spi_a_slen_hmc7044,
  output        spi_a_cs_adf4371,
  output        spi_a_csb_ad9213,
  output        spi_a_clk,
  inout         spi_a_data,
  // ADC
  output        adc_a_pdwn,
  output        adc_a_rstb,
  inout         adc_a_gpio0,
  inout         adc_a_gpio1,
  inout         adc_a_gpio2,
  inout         adc_a_gpio3,
  inout         adc_a_gpio4,
  // JESD interface
  input         jesd_a_ref_clk0_p,
  input         jesd_a_ref_clk0_n,
  input         jesd_a_ref_clk1_p,
  input         jesd_a_ref_clk1_n,
  input         jesd_a_sysref1_clk_p,
  input         jesd_a_sysref1_clk_n,
  output        jesd_a_syncinb_p,
  input [7:0]   jesd_a_serdes_0_p,
  input [7:0]   jesd_a_serdes_0_n,
  input [7:0]   jesd_a_serdes_1_p,
  input [7:0]   jesd_a_serdes_1_n,
  // Data Output Interface
  output [11:0] adc_a_dout_0,
  output [11:0] adc_a_dout_1,
  output [11:0] adc_a_dout_2,
  output [11:0] adc_a_dout_3,
  output [11:0] adc_a_dout_4,
  output [11:0] adc_a_dout_5,
  output [11:0] adc_a_dout_6,
  output [11:0] adc_a_dout_7,
  output [11:0] adc_a_dout_8,
  output [11:0] adc_a_dout_9,
  output [11:0] adc_a_dout_10,
  output [11:0] adc_a_dout_11,
  output [11:0] adc_a_dout_12,
  output [11:0] adc_a_dout_13,
  output [11:0] adc_a_dout_14,
  output [11:0] adc_a_dout_15,
  output [11:0] adc_a_dout_16,
  output [11:0] adc_a_dout_17,
  output [11:0] adc_a_dout_18,
  output [11:0] adc_a_dout_19,
  output [11:0] adc_a_dout_20,
  output [11:0] adc_a_dout_21,
  output [11:0] adc_a_dout_22,
  output [11:0] adc_a_dout_23,
  output [11:0] adc_a_dout_24,
  output [11:0] adc_a_dout_25,
  output [11:0] adc_a_dout_26,
  output [11:0] adc_a_dout_27,
  output [11:0] adc_a_dout_28,
  output [11:0] adc_a_dout_29,
  output [11:0] adc_a_dout_30,
  output [11:0] adc_a_dout_31,
  output        adc_a_clkout, // Clock domain for adc_a_dout*. (Hopefully all adc_*_dout are on the same domain)
  output [2:0]  locked_a,
  //// FMC B
  // HMC
  output        hmc_b_sync,
  output        hmc_b_reset,
  inout         hmc_b_gpio1,
  inout         hmc_b_gpio2,
  inout         hmc_b_gpio3,
  inout         hmc_b_gpio4,
  // SPI
  output        spi_b_slen_hmc7044,
  output        spi_b_cs_adf4371,
  output        spi_b_csb_ad9213,
  output        spi_b_clk,
  inout         spi_b_data,
  // ADC
  output        adc_b_pdwn,
  output        adc_b_rstb,
  inout         adc_b_gpio0,
  inout         adc_b_gpio1,
  inout         adc_b_gpio2,
  inout         adc_b_gpio3,
  inout         adc_b_gpio4,
  // JESD interface
  input         jesd_b_ref_clk0_p,
  input         jesd_b_ref_clk0_n,
  input         jesd_b_ref_clk1_p,
  input         jesd_b_ref_clk1_n,
  input         jesd_b_sysref1_clk_p,
  input         jesd_b_sysref1_clk_n,
  output        jesd_b_syncinb_p,
  input [7:0]   jesd_b_serdes_0_p,
  input [7:0]   jesd_b_serdes_0_n,
  input [7:0]   jesd_b_serdes_1_p,
  input [7:0]   jesd_b_serdes_1_n,
  // Data Output Interface
  output [11:0] adc_b_dout_0,
  output [11:0] adc_b_dout_1,
  output [11:0] adc_b_dout_2,
  output [11:0] adc_b_dout_3,
  output [11:0] adc_b_dout_4,
  output [11:0] adc_b_dout_5,
  output [11:0] adc_b_dout_6,
  output [11:0] adc_b_dout_7,
  output [11:0] adc_b_dout_8,
  output [11:0] adc_b_dout_9,
  output [11:0] adc_b_dout_10,
  output [11:0] adc_b_dout_11,
  output [11:0] adc_b_dout_12,
  output [11:0] adc_b_dout_13,
  output [11:0] adc_b_dout_14,
  output [11:0] adc_b_dout_15,
  output [11:0] adc_b_dout_16,
  output [11:0] adc_b_dout_17,
  output [11:0] adc_b_dout_18,
  output [11:0] adc_b_dout_19,
  output [11:0] adc_b_dout_20,
  output [11:0] adc_b_dout_21,
  output [11:0] adc_b_dout_22,
  output [11:0] adc_b_dout_23,
  output [11:0] adc_b_dout_24,
  output [11:0] adc_b_dout_25,
  output [11:0] adc_b_dout_26,
  output [11:0] adc_b_dout_27,
  output [11:0] adc_b_dout_28,
  output [11:0] adc_b_dout_29,
  output [11:0] adc_b_dout_30,
  output [11:0] adc_b_dout_31,
  output        adc_b_clkout, // Clock domain for adc_b_dout*. (Hopefully all adc_*_dout are on the same domain)
  output [2:0]  locked_b,
  //// FMC C
  // HMC
  output        hmc_c_sync,
  output        hmc_c_reset,
  inout         hmc_c_gpio1,
  inout         hmc_c_gpio2,
  inout         hmc_c_gpio3,
  inout         hmc_c_gpio4,
  // SPI
  output        spi_c_slen_hmc7044,
  output        spi_c_cs_adf4371,
  output        spi_c_csb_ad9213,
  output        spi_c_clk,
  inout         spi_c_data,
  // ADC
  output        adc_c_pdwn,
  output        adc_c_rstb,
  inout         adc_c_gpio0,
  inout         adc_c_gpio1,
  inout         adc_c_gpio2,
  inout         adc_c_gpio3,
  inout         adc_c_gpio4,
  // JESD interface
  input         jesd_c_ref_clk0_p,
  input         jesd_c_ref_clk0_n,
  input         jesd_c_ref_clk1_p,
  input         jesd_c_ref_clk1_n,
  input         jesd_c_sysref1_clk_p,
  input         jesd_c_sysref1_clk_n,
  output        jesd_c_syncinb_p,
  input [7:0]   jesd_c_serdes_0_p,
  input [7:0]   jesd_c_serdes_0_n,
  input [7:0]   jesd_c_serdes_1_p,
  input [7:0]   jesd_c_serdes_1_n,
  // Data Output Interface
  output [11:0] adc_c_dout_0,
  output [11:0] adc_c_dout_1,
  output [11:0] adc_c_dout_2,
  output [11:0] adc_c_dout_3,
  output [11:0] adc_c_dout_4,
  output [11:0] adc_c_dout_5,
  output [11:0] adc_c_dout_6,
  output [11:0] adc_c_dout_7,
  output [11:0] adc_c_dout_8,
  output [11:0] adc_c_dout_9,
  output [11:0] adc_c_dout_10,
  output [11:0] adc_c_dout_11,
  output [11:0] adc_c_dout_12,
  output [11:0] adc_c_dout_13,
  output [11:0] adc_c_dout_14,
  output [11:0] adc_c_dout_15,
  output [11:0] adc_c_dout_16,
  output [11:0] adc_c_dout_17,
  output [11:0] adc_c_dout_18,
  output [11:0] adc_c_dout_19,
  output [11:0] adc_c_dout_20,
  output [11:0] adc_c_dout_21,
  output [11:0] adc_c_dout_22,
  output [11:0] adc_c_dout_23,
  output [11:0] adc_c_dout_24,
  output [11:0] adc_c_dout_25,
  output [11:0] adc_c_dout_26,
  output [11:0] adc_c_dout_27,
  output [11:0] adc_c_dout_28,
  output [11:0] adc_c_dout_29,
  output [11:0] adc_c_dout_30,
  output [11:0] adc_c_dout_31,
  output        adc_c_clkout, // Clock domain for adc_c_dout*. (Hopefully all adc_*_dout are on the same domain)
  output [2:0]  locked_c,
  //// FMC D
  // HMC
  output        hmc_d_sync,
  output        hmc_d_reset,
  inout         hmc_d_gpio1,
  inout         hmc_d_gpio2,
  inout         hmc_d_gpio3,
  inout         hmc_d_gpio4,
  // SPI
  output        spi_d_slen_hmc7044,
  output        spi_d_cs_adf4371,
  output        spi_d_csb_ad9213,
  output        spi_d_clk,
  inout         spi_d_data,
  // ADC
  output        adc_d_pdwn,
  output        adc_d_rstb,
  inout         adc_d_gpio0,
  inout         adc_d_gpio1,
  inout         adc_d_gpio2,
  inout         adc_d_gpio3,
  inout         adc_d_gpio4,
  // JESD interface
  input         jesd_d_ref_clk0_p,
  input         jesd_d_ref_clk0_n,
  input         jesd_d_ref_clk1_p,
  input         jesd_d_ref_clk1_n,
  input         jesd_d_sysref1_clk_p,
  input         jesd_d_sysref1_clk_n,
  output        jesd_d_syncinb_p,
  input [7:0]   jesd_d_serdes_0_p,
  input [7:0]   jesd_d_serdes_0_n,
  input [7:0]   jesd_d_serdes_1_p,
  input [7:0]   jesd_d_serdes_1_n,
  // Data Output Interface
  output [11:0] adc_d_dout_0,
  output [11:0] adc_d_dout_1,
  output [11:0] adc_d_dout_2,
  output [11:0] adc_d_dout_3,
  output [11:0] adc_d_dout_4,
  output [11:0] adc_d_dout_5,
  output [11:0] adc_d_dout_6,
  output [11:0] adc_d_dout_7,
  output [11:0] adc_d_dout_8,
  output [11:0] adc_d_dout_9,
  output [11:0] adc_d_dout_10,
  output [11:0] adc_d_dout_11,
  output [11:0] adc_d_dout_12,
  output [11:0] adc_d_dout_13,
  output [11:0] adc_d_dout_14,
  output [11:0] adc_d_dout_15,
  output [11:0] adc_d_dout_16,
  output [11:0] adc_d_dout_17,
  output [11:0] adc_d_dout_18,
  output [11:0] adc_d_dout_19,
  output [11:0] adc_d_dout_20,
  output [11:0] adc_d_dout_21,
  output [11:0] adc_d_dout_22,
  output [11:0] adc_d_dout_23,
  output [11:0] adc_d_dout_24,
  output [11:0] adc_d_dout_25,
  output [11:0] adc_d_dout_26,
  output [11:0] adc_d_dout_27,
  output [11:0] adc_d_dout_28,
  output [11:0] adc_d_dout_29,
  output [11:0] adc_d_dout_30,
  output [11:0] adc_d_dout_31,
  output        adc_d_clkout, // Clock domain for adc_d_dout*. (Hopefully all adc_*_dout are on the same domain)
  output [2:0]  locked_d
);

wire clk_200_ibuf;
wire clk_200;

IBUFDS clk_200_ibuf_inst (
  .I(clk_200_p),
  .IB(clk_200_n),
  .O(clk_200_ibuf)
);

BUFG clk_200_bufg (
  .I(clk_200_ibuf),
  .O(clk_200)
);

generate
if (USE_FMC_A)
  ad9213_fmc_a_top ad9213_top_a_inst (
    .clk_200(clk_200),
    .reset(reset),
    .adc_clkout(adc_a_clkout),
    .uart_txd(1'b0),
    .uart_rxd(),

    .hmc_sync(hmc_a_sync),
    .hmc_reset(hmc_a_reset),
    .hmc_gpio1(hmc_a_gpio1),
    .hmc_gpio2(hmc_a_gpio2),
    .hmc_gpio3(hmc_a_gpio3),
    .hmc_gpio4(hmc_a_gpio4),

    .spi_slen_hmc7044(spi_a_slen_hmc7044),
    .spi_cs_adf4371(spi_a_cs_adf4371),
    .spi_csb_ad9213(spi_a_csb_ad9213),
    .spi_clk(spi_a_clk),
    .spi_data(spi_a_data),

    .adc_pdwn(adc_a_pdwn),
    .adc_rstb(adc_a_rstb),
    .adc_gpio0(adc_a_gpio0),
    .adc_gpio1(adc_a_gpio1),
    .adc_gpio2(adc_a_gpio2),
    .adc_gpio3(adc_a_gpio3),
    .adc_gpio4(adc_a_gpio4),

    .jesd_ref_clk0_p(jesd_a_ref_clk0_p),
    .jesd_ref_clk0_n(jesd_a_ref_clk0_n),
    .jesd_ref_clk1_p(jesd_a_ref_clk1_p),
    .jesd_ref_clk1_n(jesd_a_ref_clk1_n),
    .jesd_sysref1_clk_p(jesd_a_sysref1_clk_p),
    .jesd_sysref1_clk_n(jesd_a_sysref1_clk_n),
    .jesd_syncinb_p(jesd_a_syncinb_p),
    .serdes_0_p(jesd_a_serdes_0_p),
    .serdes_0_n(jesd_a_serdes_0_n),
    .serdes_1_p(jesd_a_serdes_1_p),
    .serdes_1_n(jesd_a_serdes_1_n),

    .adc_dout_0(adc_a_dout_0),
    .adc_dout_1(adc_a_dout_1),
    .adc_dout_2(adc_a_dout_2),
    .adc_dout_3(adc_a_dout_3),
    .adc_dout_4(adc_a_dout_4),
    .adc_dout_5(adc_a_dout_5),
    .adc_dout_6(adc_a_dout_6),
    .adc_dout_7(adc_a_dout_7),
    .adc_dout_8(adc_a_dout_8),
    .adc_dout_9(adc_a_dout_9),
    .adc_dout_10(adc_a_dout_10),
    .adc_dout_11(adc_a_dout_11),
    .adc_dout_12(adc_a_dout_12),
    .adc_dout_13(adc_a_dout_13),
    .adc_dout_14(adc_a_dout_14),
    .adc_dout_15(adc_a_dout_15),
    .adc_dout_16(adc_a_dout_16),
    .adc_dout_17(adc_a_dout_17),
    .adc_dout_18(adc_a_dout_18),
    .adc_dout_19(adc_a_dout_19),
    .adc_dout_20(adc_a_dout_20),
    .adc_dout_21(adc_a_dout_21),
    .adc_dout_22(adc_a_dout_22),
    .adc_dout_23(adc_a_dout_23),
    .adc_dout_24(adc_a_dout_24),
    .adc_dout_25(adc_a_dout_25),
    .adc_dout_26(adc_a_dout_26),
    .adc_dout_27(adc_a_dout_27),
    .adc_dout_28(adc_a_dout_28),
    .adc_dout_29(adc_a_dout_29),
    .adc_dout_30(adc_a_dout_30),
    .adc_dout_31(adc_a_dout_31),
    .locked(locked_a)
  );
endgenerate

generate
if (USE_FMC_B)
  ad9213_fmc_b_top ad9213_top_b_inst (
    .clk_200(clk_200),
    .reset(reset),
    .adc_clkout(adc_b_clkout),
    .uart_txd(1'b0),
    .uart_rxd(),

    .hmc_sync(hmc_b_sync),
    .hmc_reset(hmc_b_reset),
    .hmc_gpio1(hmc_b_gpio1),
    .hmc_gpio2(hmc_b_gpio2),
    .hmc_gpio3(hmc_b_gpio3),
    .hmc_gpio4(hmc_b_gpio4),

    .spi_slen_hmc7044(spi_b_slen_hmc7044),
    .spi_cs_adf4371(spi_b_cs_adf4371),
    .spi_csb_ad9213(spi_b_csb_ad9213),
    .spi_clk(spi_b_clk),
    .spi_data(spi_b_data),

    .adc_pdwn(adc_b_pdwn),
    .adc_rstb(adc_b_rstb),
    .adc_gpio0(adc_b_gpio0),
    .adc_gpio1(adc_b_gpio1),
    .adc_gpio2(adc_b_gpio2),
    .adc_gpio3(adc_b_gpio3),
    .adc_gpio4(adc_b_gpio4),

    .jesd_ref_clk0_p(jesd_b_ref_clk0_p),
    .jesd_ref_clk0_n(jesd_b_ref_clk0_n),
    .jesd_ref_clk1_p(jesd_b_ref_clk1_p),
    .jesd_ref_clk1_n(jesd_b_ref_clk1_n),
    .jesd_sysref1_clk_p(jesd_b_sysref1_clk_p),
    .jesd_sysref1_clk_n(jesd_b_sysref1_clk_n),
    .jesd_syncinb_p(jesd_b_syncinb_p),
    .serdes_0_p(jesd_b_serdes_0_p),
    .serdes_0_n(jesd_b_serdes_0_n),
    .serdes_1_p(jesd_b_serdes_1_p),
    .serdes_1_n(jesd_b_serdes_1_n),

    .adc_dout_0(adc_b_dout_0),
    .adc_dout_1(adc_b_dout_1),
    .adc_dout_2(adc_b_dout_2),
    .adc_dout_3(adc_b_dout_3),
    .adc_dout_4(adc_b_dout_4),
    .adc_dout_5(adc_b_dout_5),
    .adc_dout_6(adc_b_dout_6),
    .adc_dout_7(adc_b_dout_7),
    .adc_dout_8(adc_b_dout_8),
    .adc_dout_9(adc_b_dout_9),
    .adc_dout_10(adc_b_dout_10),
    .adc_dout_11(adc_b_dout_11),
    .adc_dout_12(adc_b_dout_12),
    .adc_dout_13(adc_b_dout_13),
    .adc_dout_14(adc_b_dout_14),
    .adc_dout_15(adc_b_dout_15),
    .adc_dout_16(adc_b_dout_16),
    .adc_dout_17(adc_b_dout_17),
    .adc_dout_18(adc_b_dout_18),
    .adc_dout_19(adc_b_dout_19),
    .adc_dout_20(adc_b_dout_20),
    .adc_dout_21(adc_b_dout_21),
    .adc_dout_22(adc_b_dout_22),
    .adc_dout_23(adc_b_dout_23),
    .adc_dout_24(adc_b_dout_24),
    .adc_dout_25(adc_b_dout_25),
    .adc_dout_26(adc_b_dout_26),
    .adc_dout_27(adc_b_dout_27),
    .adc_dout_28(adc_b_dout_28),
    .adc_dout_29(adc_b_dout_29),
    .adc_dout_30(adc_b_dout_30),
    .adc_dout_31(adc_b_dout_31),
    .locked(locked_b)
  );
endgenerate

generate
if (USE_FMC_C)
  ad9213_fmc_c_top ad9213_top_c_inst (
    .clk_200(clk_200),
    .reset(reset),
    .adc_clkout(adc_c_clkout),
    .uart_txd(uart_txd),
    .uart_rxd(uart_rxd),

    .hmc_sync(hmc_c_sync),
    .hmc_reset(hmc_c_reset),
    .hmc_gpio1(hmc_c_gpio1),
    .hmc_gpio2(hmc_c_gpio2),
    .hmc_gpio3(hmc_c_gpio3),
    .hmc_gpio4(hmc_c_gpio4),

    .spi_slen_hmc7044(spi_c_slen_hmc7044),
    .spi_cs_adf4371(spi_c_cs_adf4371),
    .spi_csb_ad9213(spi_c_csb_ad9213),
    .spi_clk(spi_c_clk),
    .spi_data(spi_c_data),

    .adc_pdwn(adc_c_pdwn),
    .adc_rstb(adc_c_rstb),
    .adc_gpio0(adc_c_gpio0),
    .adc_gpio1(adc_c_gpio1),
    .adc_gpio2(adc_c_gpio2),
    .adc_gpio3(adc_c_gpio3),
    .adc_gpio4(adc_c_gpio4),

    .jesd_ref_clk0_p(jesd_c_ref_clk0_p),
    .jesd_ref_clk0_n(jesd_c_ref_clk0_n),
    .jesd_ref_clk1_p(jesd_c_ref_clk1_p),
    .jesd_ref_clk1_n(jesd_c_ref_clk1_n),
    .jesd_sysref1_clk_p(jesd_c_sysref1_clk_p),
    .jesd_sysref1_clk_n(jesd_c_sysref1_clk_n),
    .jesd_syncinb_p(jesd_c_syncinb_p),
    .serdes_0_p(jesd_c_serdes_0_p),
    .serdes_0_n(jesd_c_serdes_0_n),
    .serdes_1_p(jesd_c_serdes_1_p),
    .serdes_1_n(jesd_c_serdes_1_n),

    .adc_dout_0(adc_c_dout_0),
    .adc_dout_1(adc_c_dout_1),
    .adc_dout_2(adc_c_dout_2),
    .adc_dout_3(adc_c_dout_3),
    .adc_dout_4(adc_c_dout_4),
    .adc_dout_5(adc_c_dout_5),
    .adc_dout_6(adc_c_dout_6),
    .adc_dout_7(adc_c_dout_7),
    .adc_dout_8(adc_c_dout_8),
    .adc_dout_9(adc_c_dout_9),
    .adc_dout_10(adc_c_dout_10),
    .adc_dout_11(adc_c_dout_11),
    .adc_dout_12(adc_c_dout_12),
    .adc_dout_13(adc_c_dout_13),
    .adc_dout_14(adc_c_dout_14),
    .adc_dout_15(adc_c_dout_15),
    .adc_dout_16(adc_c_dout_16),
    .adc_dout_17(adc_c_dout_17),
    .adc_dout_18(adc_c_dout_18),
    .adc_dout_19(adc_c_dout_19),
    .adc_dout_20(adc_c_dout_20),
    .adc_dout_21(adc_c_dout_21),
    .adc_dout_22(adc_c_dout_22),
    .adc_dout_23(adc_c_dout_23),
    .adc_dout_24(adc_c_dout_24),
    .adc_dout_25(adc_c_dout_25),
    .adc_dout_26(adc_c_dout_26),
    .adc_dout_27(adc_c_dout_27),
    .adc_dout_28(adc_c_dout_28),
    .adc_dout_29(adc_c_dout_29),
    .adc_dout_30(adc_c_dout_30),
    .adc_dout_31(adc_c_dout_31),
    .locked(locked_c)
  );
endgenerate

generate
if (USE_FMC_D)
  ad9213_fmc_d_top ad9213_top_d_inst (
    .clk_200(clk_200),
    .reset(reset),
    .adc_clkout(adc_d_clkout),
    .uart_txd(1'b0),
    .uart_rxd(),

    .hmc_sync(hmc_d_sync),
    .hmc_reset(hmc_d_reset),
    .hmc_gpio1(hmc_d_gpio1),
    .hmc_gpio2(hmc_d_gpio2),
    .hmc_gpio3(hmc_d_gpio3),
    .hmc_gpio4(hmc_d_gpio4),

    .spi_slen_hmc7044(spi_d_slen_hmc7044),
    .spi_cs_adf4371(spi_d_cs_adf4371),
    .spi_csb_ad9213(spi_d_csb_ad9213),
    .spi_clk(spi_d_clk),
    .spi_data(spi_d_data),

    .adc_pdwn(adc_d_pdwn),
    .adc_rstb(adc_d_rstb),
    .adc_gpio0(adc_d_gpio0),
    .adc_gpio1(adc_d_gpio1),
    .adc_gpio2(adc_d_gpio2),
    .adc_gpio3(adc_d_gpio3),
    .adc_gpio4(adc_d_gpio4),

    .jesd_ref_clk0_p(jesd_d_ref_clk0_p),
    .jesd_ref_clk0_n(jesd_d_ref_clk0_n),
    .jesd_ref_clk1_p(jesd_d_ref_clk1_p),
    .jesd_ref_clk1_n(jesd_d_ref_clk1_n),
    .jesd_sysref1_clk_p(jesd_d_sysref1_clk_p),
    .jesd_sysref1_clk_n(jesd_d_sysref1_clk_n),
    .jesd_syncinb_p(jesd_d_syncinb_p),
    .serdes_0_p(jesd_d_serdes_0_p),
    .serdes_0_n(jesd_d_serdes_0_n),
    .serdes_1_p(jesd_d_serdes_1_p),
    .serdes_1_n(jesd_d_serdes_1_n),

    .adc_dout_0(adc_d_dout_0),
    .adc_dout_1(adc_d_dout_1),
    .adc_dout_2(adc_d_dout_2),
    .adc_dout_3(adc_d_dout_3),
    .adc_dout_4(adc_d_dout_4),
    .adc_dout_5(adc_d_dout_5),
    .adc_dout_6(adc_d_dout_6),
    .adc_dout_7(adc_d_dout_7),
    .adc_dout_8(adc_d_dout_8),
    .adc_dout_9(adc_d_dout_9),
    .adc_dout_10(adc_d_dout_10),
    .adc_dout_11(adc_d_dout_11),
    .adc_dout_12(adc_d_dout_12),
    .adc_dout_13(adc_d_dout_13),
    .adc_dout_14(adc_d_dout_14),
    .adc_dout_15(adc_d_dout_15),
    .adc_dout_16(adc_d_dout_16),
    .adc_dout_17(adc_d_dout_17),
    .adc_dout_18(adc_d_dout_18),
    .adc_dout_19(adc_d_dout_19),
    .adc_dout_20(adc_d_dout_20),
    .adc_dout_21(adc_d_dout_21),
    .adc_dout_22(adc_d_dout_22),
    .adc_dout_23(adc_d_dout_23),
    .adc_dout_24(adc_d_dout_24),
    .adc_dout_25(adc_d_dout_25),
    .adc_dout_26(adc_d_dout_26),
    .adc_dout_27(adc_d_dout_27),
    .adc_dout_28(adc_d_dout_28),
    .adc_dout_29(adc_d_dout_29),
    .adc_dout_30(adc_d_dout_30),
    .adc_dout_31(adc_d_dout_31),
    .locked(locked_d)
  );
endgenerate

endmodule
