`timescale 1ns/100ps

module htg_ad9213_quad_top #(
  parameter USE_CORE_A=1,
  parameter USE_CORE_B=1,
  parameter USE_CORE_C=1,
  parameter USE_CORE_D=0
  ) (
  // 200MHz external clock
  input         clk_200_p,
  input         clk_200_n,
  // Software reset, driven from Simulink
  input         reset,
  // External UART pins
  input         uart_txd,
  output        uart_rxd,
  //// FMC A
  // HMC
  output        hmc_a_sync,
  output        hmc_a_reset,
  inout         hmc_a_gpio1,
  inout         hmc_a_gpio2,
  inout         hmc_a_gpio3,
  inout         hmc_a_gpio4,
  // SPI
  output        spi_a_slen_hmc7044,
  output        spi_a_cs_adf4371,
  output        spi_a_csb_ad9213,
  output        spi_a_clk,
  inout         spi_a_data,
  // ADC
  output        adc_a_pdwn,
  output        adc_a_rstb,
  inout         adc_a_gpio0,
  inout         adc_a_gpio1,
  inout         adc_a_gpio2,
  inout         adc_a_gpio3,
  inout         adc_a_gpio4,
  // JESD interface
  input         jesd_a_ref_clk0_p,
  input         jesd_a_ref_clk0_n,
  input         jesd_a_ref_clk1_p,
  input         jesd_a_ref_clk1_n,
  input         jesd_a_sysref1_clk_p,
  input         jesd_a_sysref1_clk_n,
  output        jesd_a_syncinb_p,
  input [7:0]   jesd_a_serdes_0_p,
  input [7:0]   jesd_a_serdes_0_n,
  input [7:0]   jesd_a_serdes_1_p,
  input [7:0]   jesd_a_serdes_1_n,
  // Data Output Interface
  output [11:0] adc_a_dout_0,
  output [11:0] adc_a_dout_1,
  output [11:0] adc_a_dout_2,
  output [11:0] adc_a_dout_3,
  output [11:0] adc_a_dout_4,
  output [11:0] adc_a_dout_5,
  output [11:0] adc_a_dout_6,
  output [11:0] adc_a_dout_7,
  output [11:0] adc_a_dout_8,
  output [11:0] adc_a_dout_9,
  output [11:0] adc_a_dout_10,
  output [11:0] adc_a_dout_11,
  output [11:0] adc_a_dout_12,
  output [11:0] adc_a_dout_13,
  output [11:0] adc_a_dout_14,
  output [11:0] adc_a_dout_15,
  output [11:0] adc_a_dout_16,
  output [11:0] adc_a_dout_17,
  output [11:0] adc_a_dout_18,
  output [11:0] adc_a_dout_19,
  output [11:0] adc_a_dout_20,
  output [11:0] adc_a_dout_21,
  output [11:0] adc_a_dout_22,
  output [11:0] adc_a_dout_23,
  output [11:0] adc_a_dout_24,
  output [11:0] adc_a_dout_25,
  output [11:0] adc_a_dout_26,
  output [11:0] adc_a_dout_27,
  output [11:0] adc_a_dout_28,
  output [11:0] adc_a_dout_29,
  output [11:0] adc_a_dout_30,
  output [11:0] adc_a_dout_31,
  output        adc_a_clkout, // Clock domain for adc_a_dout*. (Hopefully all adc_*_dout are on the same domain)
  //// FMC B
  // HMC
  output        hmc_b_sync,
  output        hmc_b_reset,
  inout         hmc_b_gpio1,
  inout         hmc_b_gpio2,
  inout         hmc_b_gpio3,
  inout         hmc_b_gpio4,
  // SPI
  output        spi_b_slen_hmc7044,
  output        spi_b_cs_adf4371,
  output        spi_b_csb_ad9213,
  output        spi_b_clk,
  inout         spi_b_data,
  // ADC
  output        adc_b_pdwn,
  output        adc_b_rstb,
  inout         adc_b_gpio0,
  inout         adc_b_gpio1,
  inout         adc_b_gpio2,
  inout         adc_b_gpio3,
  inout         adc_b_gpio4,
  // JESD interface
  input         jesd_b_ref_clk0_p,
  input         jesd_b_ref_clk0_n,
  input         jesd_b_ref_clk1_p,
  input         jesd_b_ref_clk1_n,
  input         jesd_b_sysref1_clk_p,
  input         jesd_b_sysref1_clk_n,
  output        jesd_b_syncinb_p,
  input [7:0]   jesd_b_serdes_0_p,
  input [7:0]   jesd_b_serdes_0_n,
  input [7:0]   jesd_b_serdes_1_p,
  input [7:0]   jesd_b_serdes_1_n,
  // Data Output Interface
  output [11:0] adc_b_dout_0,
  output [11:0] adc_b_dout_1,
  output [11:0] adc_b_dout_2,
  output [11:0] adc_b_dout_3,
  output [11:0] adc_b_dout_4,
  output [11:0] adc_b_dout_5,
  output [11:0] adc_b_dout_6,
  output [11:0] adc_b_dout_7,
  output [11:0] adc_b_dout_8,
  output [11:0] adc_b_dout_9,
  output [11:0] adc_b_dout_10,
  output [11:0] adc_b_dout_11,
  output [11:0] adc_b_dout_12,
  output [11:0] adc_b_dout_13,
  output [11:0] adc_b_dout_14,
  output [11:0] adc_b_dout_15,
  output [11:0] adc_b_dout_16,
  output [11:0] adc_b_dout_17,
  output [11:0] adc_b_dout_18,
  output [11:0] adc_b_dout_19,
  output [11:0] adc_b_dout_20,
  output [11:0] adc_b_dout_21,
  output [11:0] adc_b_dout_22,
  output [11:0] adc_b_dout_23,
  output [11:0] adc_b_dout_24,
  output [11:0] adc_b_dout_25,
  output [11:0] adc_b_dout_26,
  output [11:0] adc_b_dout_27,
  output [11:0] adc_b_dout_28,
  output [11:0] adc_b_dout_29,
  output [11:0] adc_b_dout_30,
  output [11:0] adc_b_dout_31,
  output        adc_b_clkout, // Clock domain for adc_b_dout*. (Hopefully all adc_*_dout are on the same domain)
  //// FMC C
  // HMC
  output        hmc_c_sync,
  output        hmc_c_reset,
  inout         hmc_c_gpio1,
  inout         hmc_c_gpio2,
  inout         hmc_c_gpio3,
  inout         hmc_c_gpio4,
  // SPI
  output        spi_c_slen_hmc7044,
  output        spi_c_cs_adf4371,
  output        spi_c_csb_ad9213,
  output        spi_c_clk,
  inout         spi_c_data,
  // ADC
  output        adc_c_pdwn,
  output        adc_c_rstb,
  inout         adc_c_gpio0,
  inout         adc_c_gpio1,
  inout         adc_c_gpio2,
  inout         adc_c_gpio3,
  inout         adc_c_gpio4,
  // JESD interface
  input         jesd_c_ref_clk0_p,
  input         jesd_c_ref_clk0_n,
  input         jesd_c_ref_clk1_p,
  input         jesd_c_ref_clk1_n,
  input         jesd_c_sysref1_clk_p,
  input         jesd_c_sysref1_clk_n,
  output        jesd_c_syncinb_p,
  input [7:0]   jesd_c_serdes_0_p,
  input [7:0]   jesd_c_serdes_0_n,
  input [7:0]   jesd_c_serdes_1_p,
  input [7:0]   jesd_c_serdes_1_n,
  // Data Output Interface
  output [11:0] adc_c_dout_0,
  output [11:0] adc_c_dout_1,
  output [11:0] adc_c_dout_2,
  output [11:0] adc_c_dout_3,
  output [11:0] adc_c_dout_4,
  output [11:0] adc_c_dout_5,
  output [11:0] adc_c_dout_6,
  output [11:0] adc_c_dout_7,
  output [11:0] adc_c_dout_8,
  output [11:0] adc_c_dout_9,
  output [11:0] adc_c_dout_10,
  output [11:0] adc_c_dout_11,
  output [11:0] adc_c_dout_12,
  output [11:0] adc_c_dout_13,
  output [11:0] adc_c_dout_14,
  output [11:0] adc_c_dout_15,
  output [11:0] adc_c_dout_16,
  output [11:0] adc_c_dout_17,
  output [11:0] adc_c_dout_18,
  output [11:0] adc_c_dout_19,
  output [11:0] adc_c_dout_20,
  output [11:0] adc_c_dout_21,
  output [11:0] adc_c_dout_22,
  output [11:0] adc_c_dout_23,
  output [11:0] adc_c_dout_24,
  output [11:0] adc_c_dout_25,
  output [11:0] adc_c_dout_26,
  output [11:0] adc_c_dout_27,
  output [11:0] adc_c_dout_28,
  output [11:0] adc_c_dout_29,
  output [11:0] adc_c_dout_30,
  output [11:0] adc_c_dout_31,
  output        adc_c_clkout, // Clock domain for adc_c_dout*. (Hopefully all adc_*_dout are on the same domain)
  //// FMC D
  // HMC
  output        hmc_d_sync,
  output        hmc_d_reset,
  inout         hmc_d_gpio1,
  inout         hmc_d_gpio2,
  inout         hmc_d_gpio3,
  inout         hmc_d_gpio4,
  // SPI
  output        spi_d_slen_hmc7044,
  output        spi_d_cs_adf4371,
  output        spi_d_csb_ad9213,
  output        spi_d_clk,
  inout         spi_d_data,
  // ADC
  output        adc_d_pdwn,
  output        adc_d_rstb,
  inout         adc_d_gpio0,
  inout         adc_d_gpio1,
  inout         adc_d_gpio2,
  inout         adc_d_gpio3,
  inout         adc_d_gpio4,
  // JESD interface
  input         jesd_d_ref_clk0_p,
  input         jesd_d_ref_clk0_n,
  input         jesd_d_ref_clk1_p,
  input         jesd_d_ref_clk1_n,
  input         jesd_d_sysref1_clk_p,
  input         jesd_d_sysref1_clk_n,
  output        jesd_d_syncinb_p,
  input [7:0]   jesd_d_serdes_0_p,
  input [7:0]   jesd_d_serdes_0_n,
  input [7:0]   jesd_d_serdes_1_p,
  input [7:0]   jesd_d_serdes_1_n,
  // Data Output Interface
  output [11:0] adc_d_dout_0,
  output [11:0] adc_d_dout_1,
  output [11:0] adc_d_dout_2,
  output [11:0] adc_d_dout_3,
  output [11:0] adc_d_dout_4,
  output [11:0] adc_d_dout_5,
  output [11:0] adc_d_dout_6,
  output [11:0] adc_d_dout_7,
  output [11:0] adc_d_dout_8,
  output [11:0] adc_d_dout_9,
  output [11:0] adc_d_dout_10,
  output [11:0] adc_d_dout_11,
  output [11:0] adc_d_dout_12,
  output [11:0] adc_d_dout_13,
  output [11:0] adc_d_dout_14,
  output [11:0] adc_d_dout_15,
  output [11:0] adc_d_dout_16,
  output [11:0] adc_d_dout_17,
  output [11:0] adc_d_dout_18,
  output [11:0] adc_d_dout_19,
  output [11:0] adc_d_dout_20,
  output [11:0] adc_d_dout_21,
  output [11:0] adc_d_dout_22,
  output [11:0] adc_d_dout_23,
  output [11:0] adc_d_dout_24,
  output [11:0] adc_d_dout_25,
  output [11:0] adc_d_dout_26,
  output [11:0] adc_d_dout_27,
  output [11:0] adc_d_dout_28,
  output [11:0] adc_d_dout_29,
  output [11:0] adc_d_dout_30,
  output [11:0] adc_d_dout_31,
  output        adc_d_clkout, // Clock domain for adc_d_dout*. (Hopefully all adc_*_dout are on the same domain)
);
